module mux8_16to1_tb;
reg[7:0] a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
reg [3:0] select;
wire[7:0] o;
mux8_16to1 m8_16to1(a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15, select, o);


initial begin
$monitor("%d a0=%b, a1=%b, a2=%b, a3=%b,a4=%b, a5=%b, a6=%b, a7=%b,a8=%b, a9=%b, a10=%b, a11=%b,a12=%b,a13=%b, a14=%b, a15=%b, select=%b, o=%b", $time,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,select,o );

a0=0;
a1=0;
a2=0;
a3=0;
a4=0;
a5=0;
a6=0;
a7=0;
a8=0;
a9=0;
a10=0;
a11=0;
a12=0;
a13=0;
a14=0;
a15=0;
select=0;


#100 a0=8'b00000000;a1=8'b10000001;a2=8'b00000010;a3=8'b10000011;a4=8'b00000111;a5=8'b11000001;a6=8'b11100010;a7=8'b10101011;a8=8'b01100000;a9=8'b11100001;a10=8'b10000010;a11=8'b10111111;a12=8'b00000000;a13=8'b10100001;a14=8'b01110010;a15=8'b10010011;select=4'b0000;
#100 a0=8'b00000000;a1=8'b10000001;a2=8'b00000010;a3=8'b10000011;a4=8'b00000111;a5=8'b11000001;a6=8'b11100010;a7=8'b10101011;a8=8'b01100000;a9=8'b11100001;a10=8'b10000010;a11=8'b10111111;a12=8'b00000000;a13=8'b10100001;a14=8'b01110010;a15=8'b10010011;select=4'b0010;
#100 a0=8'b00000000;a1=8'b10000001;a2=8'b00000010;a3=8'b10000011;a4=8'b00000111;a5=8'b11000001;a6=8'b11100010;a7=8'b10101011;a8=8'b01100000;a9=8'b11100001;a10=8'b10000010;a11=8'b10111111;a12=8'b00000000;a13=8'b10100001;a14=8'b01110010;a15=8'b10010011;select=4'b0100;
#100 a0=8'b00000000;a1=8'b10000001;a2=8'b00000010;a3=8'b10000011;a4=8'b00000111;a5=8'b11000001;a6=8'b11100010;a7=8'b10101011;a8=8'b01100000;a9=8'b11100001;a10=8'b10000010;a11=8'b10111111;a12=8'b00000000;a13=8'b10100001;a14=8'b01110010;a15=8'b10010011;select=4'b1111;


end

endmodule
